`timescale 1ns/1ns

module SM1 (
    input reset, input clock, input enable, input [31:0] dataa, input [7:0]RX,
    output reg [7:0]TX, output reg [31:0] result, output reg done, output reg [2:0]estado);


    enum integer unsigned { Idle=0, CheckSum=1, TimeOut1=2, SendBack=3, TryAlarm=4, Alarm=5, Timer=6 } fstate, reg_fstate;
    
    reg [7:0]tempo = 8'b0000_0000;
    reg [7:0]timer2 = 8'b0000_0000;
    reg [7:0]timer3 = 8'b0000_0000;

    parameter [7:0]temp = 8'b1111_1111;

    reg [7:0] firstbyte = 8'b1000_0000;
    reg [7:0] secondbyte = 8'b0000_0000;
    reg [7:0] checkdado;

    reg [7:0]SendUart_old;
    reg [7:0]result_old;
    
    reg countbyte = 0; 
    reg countSend = 0;

    reg [31:0]dataa_old;
    reg [7:0]RecevUart_old;
    
    reg [7:0] SendUart;
    reg [7:0] RecevUart;

    //reg [2:0] state = SEND_STATE;
	 reg rdy_clr;  // Limpar a entrada
	 wire rdy; //controle de leitura na uart
	 wire wr_en; // controle da escrita na uart
	 wire tx_busy;
                        //input
  	uart uart_instance(.din(SendUart), .wr_en(wr_en), .clk_50m(clock), .tx(TX), .tx_busy(tx_busy), .rx(RX), .rdy(rdy), .rdy_clr(rdy_clr), .dout(RecevUart));


    always_ff @(posedge clock or posedge reset)
    begin
        if (reset) begin
            fstate <= Idle;
        end
        else begin
            fstate <= reg_fstate;
        end
        
        
    end

    always_comb begin
        estado <= reg_fstate;
        case (fstate)
            Idle: begin
                            
                TX <= 8'bx;
                result = 8'bx;
                
                estado <= Idle; 
		        $display ("Idle");
				done <= 1'b0;
                if (dataa != dataa_old)// Se tiver algo na requis para o timer
                    reg_fstate <= Timer;
                else if (rdy)// Se tiver algo vindo da UART va para o checksum
                    reg_fstate <= CheckSum;
                else
                    reg_fstate <= Idle;
            end
            CheckSum: begin
			    $display ("CheckSum");
                checkdado <= firstbyte ^ 8'b0011_0111;

                            
                TX = 8'bx;
                result = 8'bx;
                done = 0;
                estado <= CheckSum;

                if (checkdado == secondbyte && firstbyte != 8'b0000_0000) // Se o dado estiver correto e for um dado requisitado, vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para send back
                    reg_fstate <= SendBack;
                else if (checkdado != secondbyte)// Se o dado vier "corrompido" vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para o teste de alarme
                    reg_fstate <= TryAlarm;
                else if (checkdado == secondbyte && firstbyte == 8'b0000_0000)// Se o dado estiver correto e for o alarme vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para alarme
                    reg_fstate <= Alarm;
                else
                    reg_fstate <= Idle;
            end
            TimeOut1: begin
                            
                TX = 8'bx;
                
                estado <= TimeOut1;

                $display ("TimeOut1");
                reg_fstate <= Idle;

                result <= 3'b100;// CODIGO PARA TIMEOUT NO BUFFER
				done <= 1'b1;
            end
            SendBack: begin
                TX = 8'bx;
                estado <= SendBack;

                $display ("SendBack");
                reg_fstate <= Idle;

                result <= firstbyte;// CODIGO DO DADO RECEBIDO DO ARDUINO
				done <= 1'b1;
            end
            TryAlarm: begin
                $display ("TryAlarm");
                TX = 8'bx;
                done = 0;
                result = 8'bx;
                estado <= TryAlarm;

                if (rdy)// Se ainda estiver em tempo, e receber algo na UART vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para o checksum
                    begin
                        reg_fstate <= CheckSum;
                    end
                else if (timer3 >= temp)// Caso o tempo estoure vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para o idle e grave um "bug" no buffer
                    begin
                        $display("estourou bug timer");
                        result <= 4'b1011; //CODIGO PARA BUG NO BUFFER
						done <= 1'b1;
                        reg_fstate <= Idle;
                        timer3 <= 0;
                    end
                else
                    begin
                        timer3 = timer3 + 1;
                        reg_fstate <= TryAlarm;
                    end
            end
            Alarm: begin
                $display ("Alarm");
                TX = 8'b000;
                estado = Alarm;

                if (rdy)// Se chegar algo na UART vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para o checksum
                    reg_fstate <= CheckSum;
                else if ((timer2 >= temp))// se o timer estourar vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para Idle
                    reg_fstate <= Idle;
                    timer2 <= 0;

                timer2 <= timer2 + 1;
                SendUart <= 8'b000; //CODIGO PARA CALAR A BOCA DO ALARME
                result <= 3'b111;//CODIGO PARA ALARME NO BUFFER
				done <= 1'b1;
            end
            Timer: begin
                estado = Timer;
                done = 0;
                result = 8'bx;
                $display ("Timer");
                $display ("RecevUart: %b",RecevUart);
                $display ("RecevUart: %b",RecevUart_old);
                $display ("Firstbyte: %b",firstbyte);
                $display ("secondbyte: %b",secondbyte);
                if ((tempo >= temp))// Se o tempo estourar vÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ para TimeOut (de requisiÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â§ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â£o)
                    begin
                        reg_fstate <= TimeOut1;
                        tempo = 0;
                        done <= 1'b1;
                        countSend = 0;
                    end
                else if (((rdy) & (tempo < temp)))begin

                    if (countbyte == 0)begin
                        $display("if do firstbyte = %b", countbyte);
                        firstbyte <= RecevUart;
                        countbyte = 1;
                        reg_fstate <= Timer;
                        rdy_clr <= 1'b1;
                    end
                    else if (countbyte == 1)begin
                        $display("if do secondbyte, count = %b", countbyte);
                        secondbyte <= RecevUart;
                        countbyte <= 1'b0;
                        reg_fstate <= CheckSum;
                        rdy_clr <= 1'b1;
                        countSend = 0;
                    end
                end
                // Inserting 'else' block to prevent latch inference
                else
                    begin
                        tempo = tempo + 1;
                        reg_fstate <= Timer;
                    end
				if(countSend == 0)begin
                    TX = dataa[7:0];
                    SendUart <= dataa[7:0];// CODIGO DE REQUISIÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€¦Ã‚Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¬ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡ÃƒÆ’Ã¢â‚¬Å¡Ãƒâ€šÃ‚Â¡ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã¢â‚¬Â ÃƒÂ¢Ã¢â€šÂ¬Ã¢â€žÂ¢ÃƒÆ’Ã†â€™ÃƒÂ¢Ã¢â€šÂ¬Ã‚Â ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬ÃƒÂ¢Ã¢â‚¬Å¾Ã‚Â¢ÃƒÆ’Ã†â€™Ãƒâ€ Ã¢â‚¬â„¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â‚¬Å¡Ã‚Â¬Ãƒâ€šÃ‚Â ÃƒÆ’Ã†â€™Ãƒâ€šÃ‚Â¢ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¡Ãƒâ€šÃ‚Â¬ÃƒÆ’Ã‚Â¢ÃƒÂ¢Ã¢â€šÂ¬Ã…Â¾Ãƒâ€šÃ‚Â¢O VINDA DO NIOS
                    //wr_en = 1'b1;
                    countSend = 1;
                end 
            end
            default: begin
						//fstate <= Idle;
                SendUart <= 1'bx;
                result <= 1'bx;
                //$display ("Reach undefined state");
            end
        endcase

        dataa_old = dataa;
        RecevUart_old = RecevUart;
    
    end
endmodule // SM1